library verilog;
use verilog.vl_types.all;
entity Control_Motor_vlg_vec_tst is
end Control_Motor_vlg_vec_tst;
