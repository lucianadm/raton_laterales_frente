-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 01 17:08:42 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Motor_c_ADCs IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        D : IN STD_LOGIC := '0';
        I : IN STD_LOGIC := '0';
        m : IN STD_LOGIC := '0';
        fin_cuenta : IN STD_LOGIC := '0';
        MD : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        MI : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        hab_cont : OUT STD_LOGIC
    );
END Motor_c_ADCs;

ARCHITECTURE BEHAVIOR OF Motor_c_ADCs IS
    TYPE type_fstate IS (Avanza_gDer,Izquierda_cerca,Derecha_cerca,g_Der90,g_Izq90,Avanza_gIzq);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,D,I,m,fin_cuenta)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Avanza_gDer;
            MD <= "00";
            MI <= "00";
            hab_cont <= '0';
        ELSE
            MD <= "10";
            MI <= "10";
            hab_cont <= '0';
            CASE fstate IS
                WHEN Avanza_gDer =>
                    IF (((m = '0') AND (D = '1'))) THEN
                        reg_fstate <= Derecha_cerca;
                    ELSIF ((((m = '0') AND (D = '0')) AND (I = '0'))) THEN
                        reg_fstate <= Avanza_gDer;
                    ELSIF ((((m = '0') AND (D = '0')) AND (I = '1'))) THEN
                        reg_fstate <= Izquierda_cerca;
                    ELSIF ((m = '1')) THEN
                        reg_fstate <= g_Izq90;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Avanza_gDer;
                    END IF;

                    MI <= "10";

                    hab_cont <= '0';

                    MD <= "10";
                WHEN Izquierda_cerca =>
                    IF ((I = '1')) THEN
                        reg_fstate <= Izquierda_cerca;
                    ELSIF ((I = '0')) THEN
                        reg_fstate <= Avanza_gDer;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Izquierda_cerca;
                    END IF;

                    MI <= "10";

                    hab_cont <= '0';

                    MD <= "01";
                WHEN Derecha_cerca =>
                    IF ((D = '1')) THEN
                        reg_fstate <= Derecha_cerca;
                    ELSIF ((D = '0')) THEN
                        reg_fstate <= Avanza_gDer;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Derecha_cerca;
                    END IF;

                    MI <= "01";

                    hab_cont <= '0';

                    MD <= "10";
                WHEN g_Der90 =>
                    IF ((fin_cuenta = '0')) THEN
                        reg_fstate <= g_Der90;
                    ELSIF ((fin_cuenta = '1')) THEN
                        reg_fstate <= Avanza_gDer;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= g_Der90;
                    END IF;

                    MI <= "01";

                    hab_cont <= '1';

                    MD <= "10";
                WHEN g_Izq90 =>
                    IF ((fin_cuenta = '0')) THEN
                        reg_fstate <= g_Izq90;
                    ELSIF ((fin_cuenta = '1')) THEN
                        reg_fstate <= Avanza_gIzq;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= g_Izq90;
                    END IF;

                    MI <= "10";

                    hab_cont <= '1';

                    MD <= "01";
                WHEN Avanza_gIzq =>
                    IF ((m = '1')) THEN
                        reg_fstate <= g_Der90;
                    ELSIF ((((m = '0') AND (D = '0')) AND (I = '0'))) THEN
                        reg_fstate <= Avanza_gIzq;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Avanza_gIzq;
                    END IF;

                    MI <= "10";

                    hab_cont <= '0';

                    MD <= "10";
                WHEN OTHERS => 
                    MD <= "XX";
                    MI <= "XX";
                    hab_cont <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
